//                              -*- Mode: Verilog -*-
// Filename        : alu_control_tb.v
// Description     : alu_control test bench
// Author          : Patrick
// Created On      : Fri Apr 15 15:54:38 2022
// Last Modified By: Patrick
// Last Modified On: Fri Apr 15 15:54:38 2022
// Update Count    : 0
// Status          : Unknown, Use with caution!


`timescale 1ns/1ps

//-----------------------------------------------------------------------------
// Module Declaration
//-----------------------------------------------------------------------------
module alu_control_tb (/*AUTOARG*/) ;

   //-----------------------------------------------------------------------------
   // Inputs
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Outputs
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Parameters
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Internal Registers and Wires
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Instantiations
   //-----------------------------------------------------------------------------
   alu_control duv(/*AUTOINST*/);

   //-----------------------------------------------------------------------------
   // RTL
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Assigns
   //-----------------------------------------------------------------------------
   assign clk_w_i = clk_tb_i;

endmodule // alu_control_tb

// verilog-library-flags:("-y . -y ../../rtl/verilog")
