//                              -*- Mode: Verilog -*-
// Filename        : imm_gen_tb.v
// Description     : imm gen tb
// Author          : Patrick
// Created On      : Fri Apr 15 17:22:08 2022
// Last Modified By: Patrick
// Last Modified On: Fri Apr 15 17:22:08 2022
// Update Count    : 0
// Status          : Unknown, Use with caution!

`timescale 1ns/1ps

//-----------------------------------------------------------------------------
// Module Declaration
//-----------------------------------------------------------------------------
module imm_gen_tb (/*AUTOARG*/) ;


   //-----------------------------------------------------------------------------
   // Inputs
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Outputs
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Parameters
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Internal Registers and Wires
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Instantiations
   //-----------------------------------------------------------------------------
   imm_gen duv(/*AUTOINST*/);

   //-----------------------------------------------------------------------------
   // RTL
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Assigns
   //-----------------------------------------------------------------------------

endmodule // imm_gen_tb

