//                              -*- Mode: Verilog -*-
// Filename        : registers.v
// Description     : register file for cpe cpu
// Author          : Patrick
// Created On      : Fri Apr 15 17:25:46 2022
// Last Modified By: Patrick
// Last Modified On: Fri Apr 15 17:25:46 2022
// Update Count    : 0
// Status          : Unknown, Use with caution!

//-----------------------------------------------------------------------------
// Module Declaration
//-----------------------------------------------------------------------------
module registers (/*AUTOARG*/) ;


   //-----------------------------------------------------------------------------
   // Inputs
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Outputs
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Parameters
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Internal Registers and Wires
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Instantiations
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // RTL
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Assigns
   //-----------------------------------------------------------------------------

endmodule // registers

