//                              -*- Mode: Verilog -*-
// Filename        : alu_tb.v
// Description     : test bench for the ALU module
// Author          : Patrick
// Created On      : Wed Apr 20 23:04:32 2022
// Last Modified By: Patrick
// Last Modified On: Wed Apr 20 23:04:32 2022
// Update Count    : 0
// Status          : Unknown, Use with caution!

`timescale 1ns/1ps

//-----------------------------------------------------------------------------
// Module Declaration
//-----------------------------------------------------------------------------
module alu_tb (/*AUTOARG*/) ;

   //-----------------------------------------------------------------------------
   // Inputs
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Outputs
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Parameters
   //-----------------------------------------------------------------------------
   parameter TRACE = 1;
   parameter DELAY = 1;         // TODO SET PROPER

   //-----------------------------------------------------------------------------
   // Internal Registers and Wires
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Instantiations
   //-----------------------------------------------------------------------------
   cond_branch_control duv(/*AUTOINST*/);

   //-----------------------------------------------------------------------------
   // RTL
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Assigns
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Tasks
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Tests
   //-----------------------------------------------------------------------------
   if (TRACE == 1) initial begin
      $dumpfile("cond_branch_control.vcd");
      $dumpvars;
   end

   integer errors;
   initial begin
      #DELAY;
      errors = 0;
      #DELAY;

      $display("%d ns: finished with %d errors\n", $time, errors);
   end

endmodule // alu_tb

