//                              -*- Mode: Verilog -*-
// Filename        : registers_tb.v
// Description     : register tb
// Author          : Patrick
// Created On      : Fri Apr 15 17:26:18 2022
// Last Modified By: Patrick
// Last Modified On: Fri Apr 15 17:26:18 2022
// Update Count    : 0
// Status          : Unknown, Use with caution!

`timescale 1ns/1ps

//-----------------------------------------------------------------------------
// Module Declaration
//-----------------------------------------------------------------------------
module registers_tb (/*AUTOARG*/) ;


   //-----------------------------------------------------------------------------
   // Inputs
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Outputs
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Parameters
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Internal Registers and Wires
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Instantiations
   //-----------------------------------------------------------------------------
   registers duv(/*AUTOINST*/);

   //-----------------------------------------------------------------------------
   // RTL
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Assigns
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Tests
   //-----------------------------------------------------------------------------

   if (TRACE == 1) begin
      initial begin
         $dumpfile("registers.vcd");
         $dumpvars;
      end
   end
end


endmodule // registers_tb

