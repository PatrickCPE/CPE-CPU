//                              -*- Mode: Verilog -*-
// Filename        : control_tb.v
// Description     : control generator testbench
// Author          : Patrick
// Created On      : Fri Apr 15 17:10:26 2022
// Last Modified By: Patrick
// Last Modified On: Fri Apr 15 17:10:26 2022
// Update Count    : 0
// Status          : Unknown, Use with caution!

`timescale 1ns/1ps

//-----------------------------------------------------------------------------
// Module Declaration
//-----------------------------------------------------------------------------
module control_tb (/*AUTOARG*/) ;


   //-----------------------------------------------------------------------------
   // Inputs
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Outputs
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Parameters
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Internal Registers and Wires
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Instantiations
   //-----------------------------------------------------------------------------
   control duv(/*AUTOINST*/);

   //-----------------------------------------------------------------------------
   // RTL
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Assigns
   //-----------------------------------------------------------------------------

endmodule // control_tb

