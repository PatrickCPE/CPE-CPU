//                              -*- Mode: Verilog -*-
// Filename        : cpe_cpu.v
// Description     : risk-v softcore processor implementing the RV32I spec
// Author          : Patrick
// Created On      : Fri Apr 15 15:18:58 2022
// Last Modified By: Patrick
// Last Modified On: Fri Apr 15 15:18:58 2022
// Update Count    : 0
// Status          : Unknown, Use with caution!


`timescale 1ns/1ps

//-----------------------------------------------------------------------------
// Parameters
//-----------------------------------------------------------------------------
parameter BUS_WIDTH = 32;
parameter INSTRUCTION_WIDTH = 32;

//-----------------------------------------------------------------------------
// Module Declaration
//-----------------------------------------------------------------------------
module cpe_cpu (/*AUTOARG*/ ) ;

   //-----------------------------------------------------------------------------
   // Inputs
   //-----------------------------------------------------------------------------
   input wire clk_w_i;
   input wire res_w_i_h;
   input wire [(BUS_WIDTH - 1):0]instr_w_in;

   //-----------------------------------------------------------------------------
   // Outputs
   //-----------------------------------------------------------------------------
   output wire [(BUS_WIDTH - 1):0] alu_w_o;
   output wire [(BUS_WIDTH - 1):0] reg_w_o;
   output wire [(INSTRUCTION_WIDTH - 1):0] pc_w_o;
   output wire                             mem_wr_w_o_h;
   output wire                             mem_rd_w_o_h;

   //-----------------------------------------------------------------------------
   // Internal Registers and Wires
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Instantiations
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // RTL
   //-----------------------------------------------------------------------------

   //-----------------------------------------------------------------------------
   // Assigns
   //-----------------------------------------------------------------------------

endmodule // cpe_cpu

