//                              -*- Mode: Verilog -*-
// Filename        : params.v
// Description     : global parameters to be shared throughout the cpe cpu
// Author          : Patrick
// Created On      : Fri Apr 15 15:38:50 2022
// Last Modified By: Patrick
// Last Modified On: Fri Apr 15 15:38:50 2022
// Update Count    : 0
// Status          : Unknown, Use with caution!

//-----------------------------------------------------------------------------
// Parameters
//-----------------------------------------------------------------------------
parameter BUS_WIDTH = 32;
parameter INSTRUCTION_WIDTH = 32;

endmodule // name
